    Mac OS X            	   2       8                                      ATTR      8   �   �                  �   H  com.apple.macl      �   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      q/0083;6268f891;Safari;3E7125F2-554D-41BB-B371-24DD603CFC97 