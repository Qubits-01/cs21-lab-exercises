    Mac OS X            	   2       8                                      ATTR      8   �   �                  �   H  com.apple.macl      �   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      q/0083;6268f89f;Safari;54F9A6CF-AEB3-4D68-A8CD-FC1E2F79FF95 