    Mac OS X            	   2  +     ]                                      ATTR      ]    E                    H  com.apple.macl     `   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms   !   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      bplist00�3A��r��{
                            bplist00�_]https://old-uvle.upd.edu.ph/pluginfile.php/940930/mod_folder/content/0/top.sv?forcedownload=1
                            jq/0083;6274fd65;Safari;C4D382B8-5E79-4DF1-8196-91D7BEAE9BDD 