    Mac OS X            	   2  ,     ^                                      ATTR      ^    F                    H  com.apple.macl     `   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms   "   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      bplist00�3A��pG�9
                            bplist00�_^https://old-uvle.upd.edu.ph/pluginfile.php/940930/mod_folder/content/0/dmem.sv?forcedownload=1
                            kq/0083;6274fd60;Safari;E703A566-4952-49F8-B993-849C6B403CD4 