    Mac OS X            	   2       8                                      ATTR      8   �   �                  �   H  com.apple.macl      �   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      q/0083;6274fd61;Safari;9CFFF3A2-CCAB-44AB-BC29-EC643842E9F8 