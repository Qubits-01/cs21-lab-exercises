    Mac OS X            	   2  2     d                                      ATTR      d    L                    H  com.apple.macl     `   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms   (   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      bplist00�3A��p+=
                            bplist00�_dhttps://old-uvle.upd.edu.ph/pluginfile.php/940930/mod_folder/content/0/controller.sv?forcedownload=1
                            qq/0083;6274fd60;Safari;FAABB579-33AA-44B4-9D5E-73332B44EB45 