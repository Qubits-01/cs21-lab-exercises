    Mac OS X            	   2  t     �                                      ATTR      �    �                    H  com.apple.macl     `   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms   j   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      bplist00�3A���
                            bplist00�_hhttps://old-uvle.upd.edu.ph/pluginfile.php/940929/mod_folder/content/0/imem_testbench.sv?forcedownload=1_9https://old-uvle.upd.edu.ph/mod/folder/view.php?id=466482v                            �q/0083;6268f8a0;Safari;F9003536-C38F-4579-9446-9AD30F4B26BF 