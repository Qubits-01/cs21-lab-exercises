    Mac OS X            	   2       8                                      ATTR      8   �   �                  �   H  com.apple.macl      �   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      q/0083;6268f8a0;Safari;59DA3A3C-BE68-4212-9D1D-FB0BAB906B13 