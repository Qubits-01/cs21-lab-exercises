    Mac OS X            	   2  v     �                                      ATTR      �    �                    H  com.apple.macl     `   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms   l   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      bplist00�3A��	&�
                            bplist00�_jhttps://old-uvle.upd.edu.ph/pluginfile.php/937390/mod_folder/content/0/voltin_testbench.sv?forcedownload=1_9https://old-uvle.upd.edu.ph/mod/folder/view.php?id=463320x                            �q/0083;6268f892;Safari;2F0DABC7-01D7-4FE2-B8C8-8928D1F0761E 