    Mac OS X            	   2  l     �                                      ATTR      �    �                    H  com.apple.macl     `   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms   b   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      bplist00�3A��HN
                            bplist00�_`https://old-uvle.upd.edu.ph/pluginfile.php/940929/mod_folder/content/0/aludec.sv?forcedownload=1_9https://old-uvle.upd.edu.ph/mod/folder/view.php?id=466482n                            �q/0083;6268f89e;Safari;A4EC58A0-3B68-4431-AFC5-A7350B4F74A9 