    Mac OS X            	   2       8                                      ATTR      8   �   �                  �   H  com.apple.macl      �   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      q/0083;6274fd64;Safari;1C7011A5-10B9-4EAA-ACB4-BF4B821DE4AE 