    Mac OS X            	   2       8                                      ATTR      8   �   �                  �   H  com.apple.macl      �   <  com.apple.quarantine  !��6W�I��5
#�=�                                                      q/0083;6274fd63;Safari;386C29ED-F904-4142-BE36-6FE881D2D0AA 